library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address : in std_logic_vector (11 downto 0);
        dataout : out std_logic_vector (35 downto 0)
          );
end ROM;

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0);

signal memory : memory_array:= (
       "000000000000011100000000001001100001", -- MOV A,7 
       "000000000000000100000000000101100001", -- MOV B,1 
       "000000000001010100000000000000100111", -- CALL resta 
       "000000000000001100000000000000000110", -- JMP fin 
       "000000000000000000000000001001010010", -- XOR B,A 
       "000000000000000000000000000000010111", -- PUSH B 
       "000000000000000000000000001001010010", -- XOR B,A 
       "000000000000000000000000010000100010", -- AND A,B 
       "000000000000000000000000000000001000",
       "000000000000000000000000000000011000", -- POP B 
       "000000000000000000000000000000100101", -- CMP A,0 
       "000000000000111000000000000010010110", -- JEQ suma_fin 
       "000000000000000000000000000010100011", -- SHL A 
       "000000000000010000000000000000100111", -- CALL suma 
       "000000000000000000000000001001000001", -- MOV A,B 
       "000000000000000000000000000000001000",
       "000000000000000000000000000001001000", -- RET 
       "000000000000000000000000000010000011", -- NOT A 
       "000000000000000100000000000001000100", -- INC A 
       "000000000000000000000000000000001000",
       "000000000000000000000000000001001000", -- RET 
       "000000000000000000000000000000000111", -- PUSH A 
       "000000000000000000000000001001000001", -- MOV A,B 
       "000000000001000100000000000000100111", -- CALL comp2 
       "000000000000000000000000000100010001", -- MOV B,A 
       "000000000000000000000000000000001000",
       "000000000000000000000000000000101000", -- POP A 
       "000000000000010000000000000000100111", -- CALL suma 
       "000000000000000000000000000000001000",
       "000000000000000000000000000001001000", -- RET 
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000"  -- empty
       );
begin

    dataout <= memory(to_integer(unsigned(address)));

end Behavioral;