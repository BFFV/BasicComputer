library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address : in std_logic_vector (11 downto 0);
        dataout : out std_logic_vector (35 downto 0)
          );
end ROM;

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ∗∗ 12) − 1) ) of std_logic_vector (35 downto 0);
signal memory : memory_array:= (
       "000000000000000000000000000101100001", -- a = 1 
       "000000000000000100000000010001100001", -- a = 1 
       "000000000000000000000000000101100001", -- 0 = 1 
       "000000000000000100000000010001100001", -- 0 = 1 
       "000000000000000100000000000101100001", -- b = 2 
       "000000000000001000000000010001100001", -- b = 2 
       "000000000000000100000000000101100001", -- 1 = 2 
       "000000000000001000000000010001100001", -- 1 = 2 
       "000000000000001000000000000101100001", -- c = 3 
       "000000000000001100000000010001100001", -- c = 3 
       "000000000000001000000000000101100001", -- 2 = 3 
       "000000000000001100000000010001100001", -- 2 = 3 
       "000000000000001100000000000101100001", -- d = 4 
       "000000000000010000000000010001100001", -- d = 4 
       "000000000000001100000000000101100001", -- 3 = 4 
       "000000000000010000000000010001100001", -- 3 = 4 
       "000000000000010000000000000101100001", -- e = 5 
       "000000000000010100000000010001100001", -- e = 5 
       "000000000000010000000000000101100001", -- 4 = 5 
       "000000000000010100000000010001100001", -- 4 = 5 
       "000000000000000000000000001001000001", -- MOV A,B 
       "000000000000000000000000000100010001", -- MOV B,A 
       "000000000000000000000000001001100001", -- MOV A,b 
       "000000000000110000000000000101100001", -- MOV B,Ch 
       "000000000000000000000000001001110001", -- MOV A,(a) 
       "000000000000000100000000000101110001", -- MOV B,(b) 
       "000000000000000100000000000000010001", -- MOV (b),A 
       "000000000000000000000000000001000001", -- MOV (a),B 
       "000000000000000000000000011001110001", -- MOV A,(B) 
       "000000000000000000000000010101110001", -- MOV B,(B) 
       "000000000000000000000000010000010001", -- MOV (B),A 
       "000000000000000000000000010001100001", -- MOV (B),00b 
       "000000000000000000000000010000000010", -- ADD A,B 
       "000000000000000000000000001000000010", -- ADD B,A 
       "000000000000100000000000010100000010", -- ADD A,1000b 
       "000000001111111100000000010000000010", -- ADD B,FFh 
       "000000000000001000000000010110000010", -- ADD A,(c) 
       "000000000000001100000000001110000010", -- ADD B,(d) 
       "000000000000010000000000000000000010", -- ADD (e) 
       "000000000000000000000000110110000010", -- ADD A,(B) 
       "000000000000000000000000101110000010", -- ADD B,(B) 
       "000000000000000000000000010000010010", -- SUB A,B 
       "000000000000000000000000001000010010", -- SUB B,A 
       "000000000000111100000000010100010010", -- SUB A,Fh 
       "000000000000000000000000010000010010", -- SUB B,e 
       "000000000000000000000000010110010010", -- SUB A,(a) 
       "000000000000000100000000001110010010", -- SUB B,(b) 
       "000000000000001000000000000000010010", -- SUB (c) 
       "000000000000000000000000110110010010", -- SUB A,(B) 
       "000000000000000000000000101110010010", -- SUB B,(B) 
       "000000000000000000000000010000100010", -- AND A,B 
       "000000000000000000000000001000100010", -- AND B,A 
       "000000000000000000000000010100100010", -- AND A,0 
       "000000000010000100000000010000100010", -- AND B,33d 
       "000000000000000000000000010110100010", -- AND A,(a) 
       "000000000000000100000000001110100010", -- AND B,(b) 
       "000000000000001000000000000000100010", -- AND (c) 
       "000000000000000000000000110110100010", -- AND A,(B) 
       "000000000000000000000000101110100010", -- AND B,(B) 
       "000000000000000000000000010000110010", -- OR A,B 
       "000000000000000000000000001000110010", -- OR B,A 
       "000000000000000000000000010100110010", -- OR A,e 
       "000000000001001000000000010000110010", -- OR B,12h 
       "000000000000001100000000010110110010", -- OR A,(d) 
       "000000000000010000000000001110110010", -- OR B,(e) 
       "000000000000001100000000000000110010", -- OR (d) 
       "000000000000000000000000110110110010", -- OR A,(B) 
       "000000000000000000000000101110110010", -- OR B,(B) 
       "000000000000000000000000010001010010", -- XOR A,B 
       "000000000000000000000000001001010010", -- XOR B,A 
       "000000000000111100000000010101010010", -- XOR A,1111b 
       "000001000101011100000000010001010010", -- XOR B,1111d 
       "000000000000001000000000010111010010", -- XOR A,(c) 
       "000000000000001100000000001111010010", -- XOR B,(d) 
       "000000000000000000000000000001010010", -- XOR (a) 
       "000000000000000000000000110111010010", -- XOR A,(B) 
       "000000000000000000000000101111010010", -- XOR B,(B) 
       "000000000000000000000000000010000011", -- NOT A 
       "000000000000000000000000000001000011", -- NOT B,A 
       "000000000000001000000000000000000011", -- NOT (c),A 
       "000000000000000000000000000100000011", -- NOT (B),A 
       "000000000000000000000000000010100011", -- SHL A 
       "000000000000000000000000000001100011", -- SHL B,A 
       "000000000000000000000000000000100011", -- SHL (a),A 
       "000000000000000000000000000100100011", -- SHL (B),A 
       "000000000000000000000000000010110011", -- SHR A 
       "000000000000000000000000000001110011", -- SHR B,A 
       "000000000000001000000000000000110011", -- SHR (c),A 
       "000000000000000000000000000100110011", -- SHR (B),A 
       "000000000000000100000000000001000100", -- INC A 
       "000000000000000100000000000000000100", -- INC B 
       "000000000000001100000000000001100100", -- INC (d) 
       "000000000000000100000000000011100100", -- INC (B) 
       "000000000000000100000000000001010100", -- DEC A 
       "000000000000000000000000000000000101", -- CMP A,B 
       "000000000000000000000000000000100101", -- CMP A,a 
       "000000000000000000000000000000110101", -- CMP A,(a) 
       "000000000000000000000000000001110101", -- CMP A,(B) 
       "000000000101111000000000000000000110", -- JMP jump 
       "000000000101111000000000000010010110", -- JEQ jump 
       "000000000101111000000000000000010110", -- JNE jump 
       "000000000101111000000000000000110110", -- JGT jump 
       "000000000101111000000000000000100110", -- JGE jump 
       "000000000101111000000000000010100110", -- JLT jump 
       "000000000101111000000000000010110110", -- JLE jump 
       "000000000101111000000000000011000110", -- JCR jump 
       "000000000000000000000000000000000111", -- PUSH A 
       "000000000000000000000000000000010111", -- PUSH B 
       "000000000110111000000000000000100111", -- CALL none 
       "000000000111010000000000000000000110", -- JMP xd 
       "000000000000000000000000000000000000", -- NOP 
       "000000000000000000000000000000000000", -- NOP 
       "000000000000000000000000000000000000", -- NOP 
       "000000000000000000000000000000000000", -- NOP 
       "000000000000000000000000000000001000",
       "000000000000000000000000000001001000", -- RET 
       "000000000000000000000000000000001000",
       "000000000000000000000000000000101000", -- POP A 
       "000000000000000000000000000000001000",
       "000000000000000000000000000000011000", -- POP B 
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       );
begin

    dataout <= memory(to_integer(unsigned(address)));

end Behavioral;