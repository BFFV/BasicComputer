library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (
	"000000000000000000000000000101100001", -- MOV B,0
	"000000000000000000000000000001000001", -- MOV (0),B
	"000000000000001000000000000101100001", -- MOV B,2          *** Num1
	"000000000000000100000000000001000001", -- MOV (1),B
	"000000000000100100000000000101100001", -- MOV B,9          *** Num2
	"000000000000001000000000000001000001", -- MOV (2),B
	"000000000000000000000000000101100001", -- MOV B,0
	"000000000000000100000000001001110001", -- MOV A,(1)
	"000000000000001000000000000101110001", -- MOV B,(2)
	"000000000000000000000000000000100101", -- CMP A,0
	"000000000001000100000000000010010110", -- JEQ 17
	"000000000000000000000000001001110001", -- MOV A,(0)
	"000000000000000000000000000000000010", -- ADD (0)
	"000000000000000100000000001001110001", -- MOV A,(1)
	"000000000000000100000000000001010100", -- DEC A
	"000000000000000100000000000000010001", -- MOV (1),A
	"000000000000100100000000000000000110", -- JMP 9
	"000000000000000000000000001001110001", -- MOV A,(0)
	"000000000001001000000000000000000110", -- JMP 18
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000"
        ); 
begin

   dataout <= memory(to_integer(unsigned(address))); 

end Behavioral; 
