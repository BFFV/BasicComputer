library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address : in std_logic_vector (11 downto 0);
        dataout : out std_logic_vector (35 downto 0)
          );
end ROM;

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0);

signal memory : memory_array:= (
       "000000000000000000000000000101100001", -- var = 10 
       "000000000000101000000000010001100001", -- var = 10 
       "000000000000010000000000000000000110", -- JMP paso1 
       "000000000001000000000000001001100001", -- MOV A,16 
       "000000000000001100000000001001100001", -- MOV A,3 
       "000000000000010000000000000000100101", -- CMP A,4 
       "000000000000100000000000000000010110", -- JNE paso2 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000001100000000001001100001", -- MOV A,3 
       "000000000000001100000000000000100101", -- CMP A,3 
       "000000000000110000000000000010010110", -- JEQ paso3 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000101000000000001001100001", -- MOV A,10 
       "000000000000010000000000000000100101", -- CMP A,4 
       "000000000001000000000000000000110110", -- JGT paso4 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000001010000000000000000100101", -- CMP A,20 
       "000000000001001100000000000010100110", -- JLT paso5 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000100000000000000000100101", -- CMP A,8 
       "000000000001011000000000000000100110", -- JGE next1 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000000000000000000000110101", -- CMP A,(var) 
       "000000000001100100000000000000100110", -- JGE paso6 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000101100000000000000100101", -- CMP A,11 
       "000000000001110000000000000010110110", -- JLE next2 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000000000000000000000110101", -- CMP A,(var) 
       "000000000001111100000000000010110110", -- JLE paso7 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000001111111100000000001001100001", -- MOV A,255 
       "000000000000101000000000010100000010", -- ADD A,10 
       "000000000000000000000000000000000101", -- CMP A,B 
       "000000000010011100000000000011000110", -- JCR fin 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000000111100000000001001100001", -- MOV A,15 
       "000000000000111100000000000101100001", -- MOV B,15 
       "000000000010010000000000000000000110", -- JMP loop 
       "000000000001000000000000001001100001", -- MOV A,16 
       "000000000001000000000000000101100001", -- MOV B,16 
       "000000000010011100000000000000000110", -- JMP fin 
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000"  -- empty
       );
begin

    dataout <= memory(to_integer(unsigned(address)));

end Behavioral;