library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address : in std_logic_vector (11 downto 0);
        dataout : out std_logic_vector (35 downto 0)
          );
end ROM;

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0);

signal memory : memory_array:= (
       "000000000000000000000000000101100001", -- odd = 0 
       "000000000000000000000000010001100001", -- odd = 0 
       "000000000000000100000000000101100001", -- last = 0 
       "000000000000000000000000010001100001", -- last = 0 
       "000000000000001000000000000000101001", -- IN A,2 
       "000000000000000100000000010100100010", -- AND A,1 
       "000000000000000000000000000000010001", -- MOV (odd),A 
       "000000000000000000000000000000011001", -- IN B,0 
       "000000000000000000000000001001100001", -- MOV A,0 
       "000000000000000000000000000010000011", -- NOT A 
       "000000000000000000000000010110000010", -- ADD A,(odd) 
       "000000000000000000000000010001010010", -- XOR A,B 
       "000000000000000100000000000000101010", -- OUT A,1 
       "000000000000000100000000001001110001", -- MOV A,(last) 
       "000000000000000000000000000000110101", -- CMP A,(odd) 
       "000000000000010000000000000010010110", -- JEQ loop 
       "000000000000000100000000000101100001", -- MOV B,1 
       "000000000000000100000000000001010010", -- XOR (last) 
       "000000000000000100000000000000101001", -- IN A,1 
       "000000000000000000000000000000101010", -- OUT A,0 
       "000000000000010000000000000000000110", -- JMP loop 
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000"  -- empty
       );
begin

    dataout <= memory(to_integer(unsigned(address)));

end Behavioral;