library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address : in std_logic_vector (11 downto 0);
        dataout : out std_logic_vector (35 downto 0)
          );
end ROM;

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ∗∗ 12) − 1) ) of std_logic_vector (35 downto 0);
signal memory : memory_array:= (
       "000000000000000000000000000101100001", -- a = 1 
       "000000000000000100000000010001100001", -- a = 1 
       "000000000000000000000000000101100001", -- 0 = 1 
       "000000000000000100000000010001100001", -- 0 = 1 
       "000000000000000100000000000101100001", -- b = 1 
       "000000000000000100000000010001100001", -- b = 1 
       "000000000000000100000000000101100001", -- 1 = 1 
       "000000000000000100000000010001100001", -- 1 = 1 
       "000000000000001000000000000101100001", -- c = 2 
       "000000000000001000000000010001100001", -- c = 2 
       "000000000000001000000000000101100001", -- 2 = 2 
       "000000000000001000000000010001100001", -- 2 = 2 
       "000000000000001100000000000101100001", -- d = 4 
       "000000000000010000000000010001100001", -- d = 4 
       "000000000000001100000000000101100001", -- 3 = 4 
       "000000000000010000000000010001100001", -- 3 = 4 
       "000000000000000000000000001001100001", -- MOV A,0 
       "000000000000001000000000000101100001", -- MOV B,2 
       "000000000000000000000000000000000101", -- CMP A,B 
       "000000000001010000000000000010010110", -- JEQ primer_salto 
       "000000000000000100000000001001100001", -- MOV A,1 
       "000000000000000000000000010000100010", -- AND A,B 
       "000000000000000000000000000000000101", -- CMP A,B 
       "000000000001100000000000000000010110", -- JNE segundo_salto 
       "000000000000000000000000010001010010", -- XOR A,B 
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       "000000000000000000000000000000000000", -- empty
       );
begin

    dataout <= memory(to_integer(unsigned(address)));

end Behavioral;